<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.25,-1.3009,126.275,-59.7076</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>40.5,-18</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_NAND2</type>
<position>40.5,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>28.5,-17</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>28.5,-26</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>53.5,-18</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>53.5,-25</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>41,-10.5</position>
<gparam>LABEL_TEXT SR Latch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>28.5,-14.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>28.5,-23.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>53.5,-15.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>112,-18.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>112,-25.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>125,-18.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>125,-25.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>100,-15.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>100,-25</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>125,-16</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>98.5,-9</position>
<gparam>LABEL_TEXT Gated D Latch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>BA_NAND2</type>
<position>95.5,-17.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>95.5,-26.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>87,-21.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>87,-19</position>
<gparam>LABEL_TEXT W</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>79.5,-16.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_SMALL_INVERTER</type>
<position>82.5,-23.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>79.5,-14</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AE_DFF_LOW</type>
<position>44.5,-45.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUTINV_0</ID>15 </output>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clock</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>28,-43.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>BB_CLOCK</type>
<position>28.5,-50</position>
<output>
<ID>CLK</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>28,-41.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>28,-47</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>55,-43.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>55,-47.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>55,-41</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>55,-45.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>43.5,-38</position>
<gparam>LABEL_TEXT D Flip Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-18,52.5,-18</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>45.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-20.5,45.5,-18</points>
<intersection>-20.5 5</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>34.5,-20.5,45.5,-20.5</points>
<intersection>34.5 6</intersection>
<intersection>45.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>34.5,-24,34.5,-20.5</points>
<intersection>-24 7</intersection>
<intersection>-20.5 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>34.5,-24,37.5,-24</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>34.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-25,45,-22</points>
<intersection>-25 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-25,52.5,-25</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-22,45,-22</points>
<intersection>36 3</intersection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-22,36,-19</points>
<intersection>-22 2</intersection>
<intersection>-19 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-19,37.5,-19</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-17,37.5,-17</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-26,37.5,-26</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-26,37.5,-26</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-18.5,124,-18.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>117 4</intersection>
<intersection>124 14</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117,-21,117,-18.5</points>
<intersection>-21 5</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>106,-21,117,-21</points>
<intersection>106 6</intersection>
<intersection>117 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>106,-24.5,106,-21</points>
<intersection>-24.5 7</intersection>
<intersection>-21 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>106,-24.5,109,-24.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>106 6</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>124,-18.5,124,-18.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-25.5,116.5,-22.5</points>
<intersection>-25.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-25.5,124,-25.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-22.5,116.5,-22.5</points>
<intersection>107.5 3</intersection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107.5,-22.5,107.5,-19.5</points>
<intersection>-22.5 2</intersection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>107.5,-19.5,109,-19.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>107.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98.5,-17.5,109,-17.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98.5,-26.5,109,-26.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-25.5,91,-18.5</points>
<intersection>-25.5 2</intersection>
<intersection>-21.5 3</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-18.5,92.5,-18.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-25.5,92.5,-25.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89,-21.5,91,-21.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-16.5,92.5,-16.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>82.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-21.5,82.5,-16.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-27.5,82.5,-25.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-27.5,92.5,-27.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-43.5,54,-43.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-47.5,50.5,-46.5</points>
<intersection>-47.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-47.5,54,-47.5</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-46.5,50.5,-46.5</points>
<connection>
<GID>38</GID>
<name>OUTINV_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-50,37,-46.5</points>
<intersection>-50 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-46.5,41.5,-46.5</points>
<connection>
<GID>38</GID>
<name>clock</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-50,37,-50</points>
<connection>
<GID>46</GID>
<name>CLK</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-43.5,41.5,-43.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>