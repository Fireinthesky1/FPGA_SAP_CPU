james@FIRE.15140:1701069165