library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity three_ones is

end three_ones;

architecture my_arch of three_ones is

end my_arch;
