james@DESKTOP-CL1GNN2.10028:1697086000