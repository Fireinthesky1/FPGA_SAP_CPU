<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>18.6852,-9.23354,149.19,-77.275</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>55,-60.5</position>
<gparam>LABEL_TEXT c2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>87.5,-37.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>49,-58.5</position>
<gparam>LABEL_TEXT c3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_OR2</type>
<position>101,-38</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>97.5,-61</position>
<gparam>LABEL_TEXT c0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR3</type>
<position>110.5,-54.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>100,-55</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_OR2</type>
<position>88.5,-66</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AI_XOR3</type>
<position>67,-55.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>53.5,-55</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>15 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>47.5,-55</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR3</type>
<position>51.5,-68.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>44,-38</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR2</type>
<position>58,-38</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>102,-17</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>86.5,-16.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>123,-45</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>86.5,-13.5</position>
<gparam>LABEL_TEXT a0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>102,-14</position>
<gparam>LABEL_TEXT b0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>123,-42.5</position>
<gparam>LABEL_TEXT carry in</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>104,-40</position>
<gparam>LABEL_TEXT p0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>90.5,-40</position>
<gparam>LABEL_TEXT g0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>81.5,-61</position>
<gparam>LABEL_TEXT c1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>59,-17.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>43.5,-17.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>43.5,-14.5</position>
<gparam>LABEL_TEXT a1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>59,-14.5</position>
<gparam>LABEL_TEXT b1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>110.5,-76</position>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>67,-76</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>51.5,-76</position>
<input>
<ID>N_in3</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>113.5,-58.5</position>
<gparam>LABEL_TEXT sum0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>70,-60</position>
<gparam>LABEL_TEXT sum1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>56,-72.5</position>
<gparam>LABEL_TEXT carry out</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>61,-41</position>
<gparam>LABEL_TEXT p1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>46,-41.5</position>
<gparam>LABEL_TEXT g1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>82,-10</position>
<gparam>LABEL_TEXT Eight Bit Carry Lookahead Adder (work in progress)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-75,51.5,-71.5</points>
<connection>
<GID>30</GID>
<name>N_in3</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-51.5,110.5,-27</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>88.5,-27,110.5,-27</points>
<intersection>88.5 5</intersection>
<intersection>102 9</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>88.5,-34.5,88.5,-27</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-27 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>102,-35,102,-19</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-27 4</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-34.5,86.5,-18.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-29.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>86.5,-29.5,108.5,-29.5</points>
<intersection>86.5 0</intersection>
<intersection>100 8</intersection>
<intersection>108.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>108.5,-51.5,108.5,-29.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>-29.5 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>100,-35,100,-29.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-29.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-75,110.5,-57.5</points>
<connection>
<GID>28</GID>
<name>N_in3</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-52,101,-41</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-43 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53.5,-43,101,-43</points>
<intersection>53.5 5</intersection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53.5,-52,53.5,-43</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-43 4</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-63,89.5,-60</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-60 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100,-60,100,-58</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-60,100,-60</points>
<intersection>89.5 0</intersection>
<intersection>100 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-63,87.5,-40.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-47,87.5,-47</points>
<intersection>46.5 2</intersection>
<intersection>87.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>46.5,-52,46.5,-47</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-47 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-52.5,69,-51</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-70,83,-51</points>
<intersection>-70 3</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-51,83,-51</points>
<intersection>69 0</intersection>
<intersection>83 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83,-70,88.5,-70</points>
<intersection>83 1</intersection>
<intersection>88.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>88.5,-70,88.5,-69</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>-70 3</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-51.5,112.5,-45</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-45,121,-45</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>55.5 5</intersection>
<intersection>99 3</intersection>
<intersection>112.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>99,-52,99,-45</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-45 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>55.5,-52,55.5,-45</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-65.5,53.5,-58</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-61.5,47.5,-58</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>-61.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-61.5,51.5,-61.5</points>
<intersection>47.5 0</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-65.5,51.5,-61.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-61.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-65.5,44,-41</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>-65.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>44,-65.5,49.5,-65.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-35,59,-19.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-27,67,-27</points>
<intersection>45 7</intersection>
<intersection>59 0</intersection>
<intersection>67 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>45,-35,45,-27</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-27 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>67,-52.5,67,-27</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>-27 4</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-52.5,65,-29.5</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>-29.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-29.5,65,-29.5</points>
<intersection>43.5 5</intersection>
<intersection>57 18</intersection>
<intersection>65 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-35,43.5,-19.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-35 19</intersection>
<intersection>-29.5 4</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>57,-35,57,-29.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-29.5 4</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>43,-35,43.5,-35</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>43.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-52,51.5,-42</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>-42 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58,-42,58,-41</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-42,58,-42</points>
<intersection>48.5 4</intersection>
<intersection>51.5 0</intersection>
<intersection>58 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-52,48.5,-42</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-75,67,-58.5</points>
<connection>
<GID>29</GID>
<name>N_in3</name></connection>
<connection>
<GID>9</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>