module not
(
  input [bits-1:0] x_i,
  output           f_o
);

wire f_w;
nand(f_w, );

endmodule