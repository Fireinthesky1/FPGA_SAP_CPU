<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-10.7161,6.76646,99.8411,-50.875</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>66,-19</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>59,-19</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>52,-19</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>74,-1.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>70,-1.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>74,0.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>70,0.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR3</type>
<position>58,-32</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR3</type>
<position>74,-19.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>FF_GND</type>
<position>76,-14</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>82.5,-14</position>
<gparam>LABEL_TEXT Disconnected</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>FF_GND</type>
<position>60,-14</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>FF_GND</type>
<position>53,-14</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>17.5,-17.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>10.5,-17.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>3.5,-17.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>25.5,-0.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>20,-0.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>25.5,2</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>20,2</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR3</type>
<position>9.5,-30.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR3</type>
<position>25.5,-18</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>74,-42.5</position>
<input>
<ID>N_in3</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>58,-37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Carry In</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>33.5,-12</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Carry In</lparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>70.5,-42.5</position>
<input>
<ID>N_in2</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>66.5,-42.5</position>
<input>
<ID>N_in2</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>48,6</position>
<gparam>LABEL_TEXT Two Bit Ripple Carry Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-16.5,76,-15</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-16.5,74,-3.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-16.5 8</intersection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>58,-12.5,74,-12.5</points>
<intersection>58 7</intersection>
<intersection>67 5</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>67,-16,67,-12.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-12.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>58,-16,58,-12.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>74,-16.5,74,-16.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-16.5,72,-10</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>-10 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-10,70,-3.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51,-10,72,-10</points>
<intersection>51 9</intersection>
<intersection>65 4</intersection>
<intersection>70 1</intersection>
<intersection>72 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>65,-16,65,-10</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-10 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>51,-16,51,-10</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-10 2</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-16,60,-15</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-16,53,-15</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-29,60,-25.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66,-25.5,66,-22</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-25.5,66,-25.5</points>
<intersection>60 0</intersection>
<intersection>66 1</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-29,58,-25.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59,-25.5,59,-22</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,-25.5,59,-25.5</points>
<intersection>58 0</intersection>
<intersection>59 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-29,56,-25.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,-25.5,52,-22</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,-25.5,56,-25.5</points>
<intersection>52 1</intersection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-15,25.5,-2.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-11 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9.5,-11,25.5,-11</points>
<intersection>9.5 7</intersection>
<intersection>18.5 5</intersection>
<intersection>25.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>18.5,-14.5,18.5,-11</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-11 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>9.5,-14.5,9.5,-11</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-11 4</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-15,23.5,-8.5</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20,-8.5,20,-2.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-8.5,23.5,-8.5</points>
<intersection>2.5 6</intersection>
<intersection>16.5 4</intersection>
<intersection>20 1</intersection>
<intersection>23.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16.5,-14.5,16.5,-8.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>2.5,-14.5,2.5,-8.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-8.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-27.5,11.5,-24</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17.5,-24,17.5,-20.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-24,17.5,-24</points>
<intersection>11.5 0</intersection>
<intersection>17.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-27.5,9.5,-24</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-24,10.5,-20.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-24,10.5,-24</points>
<intersection>9.5 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-27.5,7.5,-24</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3.5,-24,3.5,-20.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-24,7.5,-24</points>
<intersection>3.5 1</intersection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-41.5,74,-22.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-35.5,58,-35</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-15,27.5,-12</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-12,31.5,-12</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>4.5 5</intersection>
<intersection>11.5 3</intersection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>11.5,-14.5,11.5,-12</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>4.5,-14.5,4.5,-12</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-50.5,25.5,-21</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70.5,-50.5,70.5,-43.5</points>
<connection>
<GID>43</GID>
<name>N_in2</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-50.5,70.5,-50.5</points>
<intersection>25.5 0</intersection>
<intersection>70.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-48.5,66.5,-43.5</points>
<connection>
<GID>45</GID>
<name>N_in2</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9.5,-48.5,9.5,-33.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-48.5,66.5,-48.5</points>
<intersection>9.5 1</intersection>
<intersection>66.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>