<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-6,0,171.8,-92.7</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>6.5,-15.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>6.5,-17.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>4.5,-15</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>4.5,-17.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AI_XOR2</type>
<position>23,-16.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>23,-22.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>43,-22.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>33,-22.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>43,-20</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>33,-20</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>26.5,-10.5</position>
<gparam>LABEL_TEXT half adder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>98,-13.5</position>
<gparam>LABEL_TEXT full adder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>77,-19</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>77,-21</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>75,-18.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>75,-21</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>77,-23</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>72.5,-23</position>
<gparam>LABEL_TEXT carry in</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR3</type>
<position>92.5,-21</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>10 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>92,-28</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>92,-34</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>92,-40</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>117,-34</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>125,-34</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>117,-31.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>125,-31.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_OR3</type>
<position>108,-34</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-17.5,20,-17.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-23.5,13,-17.5</points>
<intersection>-23.5 4</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13,-23.5,20,-23.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>13 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-15.5,20,-15.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-21.5,15.5,-15.5</points>
<intersection>-21.5 4</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-21.5,20,-21.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-22.5,32,-22.5</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-22.5,38,-16.5</points>
<intersection>-22.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-22.5,42,-22.5</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-16.5,38,-16.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-19,89.5,-19</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>87 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>87,-33,87,-19</points>
<intersection>-33 16</intersection>
<intersection>-27 14</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>87,-27,89,-27</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>87 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>87,-33,89,-33</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>87 13</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-23,89.5,-23</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>83 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>83,-41,83,-23</points>
<intersection>-41 14</intersection>
<intersection>-35 12</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>83,-35,89,-35</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>83 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>83,-41,89,-41</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>83 11</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-21,89.5,-21</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>85 3</intersection>
<intersection>89.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-39,85,-21</points>
<intersection>-39 6</intersection>
<intersection>-29 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>85,-29,89,-29</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>85 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>85,-39,89,-39</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>85 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>89.5,-21,89.5,-21</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-34,121,-21</points>
<intersection>-34 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-34,124,-34</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-21,121,-21</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,-34,105,-34</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-32,100,-28</points>
<intersection>-32 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-32,105,-32</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95,-28,100,-28</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-40,100,-36</points>
<intersection>-40 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-36,105,-36</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95,-40,100,-40</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-34,116,-34</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>52</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-92.7</PageViewport></page 9></circuit>