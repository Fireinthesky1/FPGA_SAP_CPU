<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-73.1163,31.7665,73.6913,-44.775</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>4.5,2.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_OR2</type>
<position>18,2</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR3</type>
<position>27.5,-14.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>17,-15</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>5.5,-26</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AI_XOR3</type>
<position>-16,-15.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND3</type>
<position>-29.5,-15</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>15 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>-35.5,-15</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR3</type>
<position>-31.5,-28.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>-39,2</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>-25,2</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>16,23.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>3.5,23.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>40,-5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>3.5,26.5</position>
<gparam>LABEL_TEXT a0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>16,26.5</position>
<gparam>LABEL_TEXT b0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>40,-2.5</position>
<gparam>LABEL_TEXT cin0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>21,0</position>
<gparam>LABEL_TEXT p0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>7.5,0</position>
<gparam>LABEL_TEXT g0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>2,-31.5</position>
<gparam>LABEL_TEXT cout0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-10,-12</position>
<gparam>LABEL_TEXT cin1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>11,23.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-1.5,23.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-1.5,26.5</position>
<gparam>LABEL_TEXT a1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>11,26.5</position>
<gparam>LABEL_TEXT b1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>-11.5,-43.5</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>-16,-43.5</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>-20.5,-43.5</position>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>31,-18.5</position>
<gparam>LABEL_TEXT sum0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-12.5,-20</position>
<gparam>LABEL_TEXT sum1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>-27.5,-32.5</position>
<gparam>LABEL_TEXT cout1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-21.5,-1</position>
<gparam>LABEL_TEXT p1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>-37,-1.5</position>
<gparam>LABEL_TEXT g1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>7.5,31</position>
<gparam>LABEL_TEXT Two Bit Carry Lookahead Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-11.5,27.5,13</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5.5,13,27.5,13</points>
<intersection>5.5 5</intersection>
<intersection>16 9</intersection>
<intersection>19 14</intersection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>5.5,5.5,5.5,13</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>13 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>16,13,16,21.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>13 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>19,5,19,13</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,5.5,3.5,21.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>10.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>3.5,10.5,25.5,10.5</points>
<intersection>3.5 0</intersection>
<intersection>17 8</intersection>
<intersection>25.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>25.5,-11.5,25.5,10.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>10.5 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>17,5,17,10.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>10.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-12,18,-1</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-3 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-29.5,-3,18,-3</points>
<intersection>-29.5 5</intersection>
<intersection>18 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-29.5,-12,-29.5,-3</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-3 4</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-23,6.5,-20</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,-20,17,-18</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-20,17,-20</points>
<intersection>6.5 0</intersection>
<intersection>17 1</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-23,4.5,-0.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-7,4.5,-7</points>
<intersection>-36.5 2</intersection>
<intersection>4.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-36.5,-12,-36.5,-7</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-12.5,-14,-11</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>0,-30,0,-11</points>
<intersection>-30 3</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-11,0,-11</points>
<intersection>-14 0</intersection>
<intersection>0 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>0,-30,5.5,-30</points>
<intersection>0 1</intersection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-30,5.5,-29</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>-30 3</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-11.5,29.5,-5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-5,38,-5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 5</intersection>
<intersection>16 3</intersection>
<intersection>29.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-12,16,-5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-27.5,-12,-27.5,-5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-25.5,-29.5,-18</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-21.5,-35.5,-18</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-35.5,-21.5,-31.5,-21.5</points>
<intersection>-35.5 0</intersection>
<intersection>-31.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-31.5,-25.5,-31.5,-21.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-21.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-25.5,-39,-1</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-25.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-39,-25.5,-33.5,-25.5</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,9,11,21.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-38,9,11,9</points>
<intersection>-38 7</intersection>
<intersection>-24 5</intersection>
<intersection>-16 9</intersection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-24,5,-24,9</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>9 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-38,5,-38,9</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>9 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-16,-12.5,-16,9</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>9 4</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-12.5,-18,10.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>10.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-40,10.5,-1.5,10.5</points>
<intersection>-40 5</intersection>
<intersection>-26 11</intersection>
<intersection>-18 0</intersection>
<intersection>-1.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-40,5,-40,10.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>10.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-1.5,10.5,-1.5,21.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>10.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-26,5,-26,10.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>10.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-12,-31.5,-2</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>-2 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-25,-2,-25,-1</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-2,-25,-2</points>
<intersection>-34.5 4</intersection>
<intersection>-31.5 0</intersection>
<intersection>-25 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-34.5,-12,-34.5,-2</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-2 2</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-42.5,-11.5,-40.5</points>
<connection>
<GID>37</GID>
<name>N_in3</name></connection>
<intersection>-40.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27.5,-40.5,27.5,-17.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-40.5,27.5,-40.5</points>
<intersection>-11.5 0</intersection>
<intersection>27.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-42.5,-16,-18.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-42.5,-20.5,-37</points>
<connection>
<GID>39</GID>
<name>N_in3</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-31.5,-37,-31.5,-31.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-31.5,-37,-20.5,-37</points>
<intersection>-31.5 1</intersection>
<intersection>-20.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 1>
<page 2>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,3.48214e-006,177.8,-92.7</PageViewport></page 9></circuit>