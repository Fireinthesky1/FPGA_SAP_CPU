$date
  Sat Nov 11 18:26:34 2023
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module tb $end
$var reg 1 ! clk $end
$var reg 1 " btn $end
$var reg 1 # rst $end
$var reg 3 $ cnt[2:0] $end
$scope module threebitcounter $end
$var reg 1 % clk $end
$var reg 1 & btn $end
$var reg 1 ' rst $end
$var reg 3 ( cnt[2:0] $end
$var reg 1 ) q0_int $end
$var reg 1 * q1_int $end
$var reg 1 + q2_int $end
$var reg 1 , btn_db $end
$scope module debouncer $end
$var reg 1 - reset $end
$var reg 1 . clk $end
$var reg 1 / sw $end
$var reg 1 0 db $end
$var reg 20 1 ctr_reg[19:0] $end
$var reg 20 2 ctr_nxt[19:0] $end
$var reg 1 3 m_tick $end
$comment state_reg is not handled $end
$comment state_nxt is not handled $end
$upscope $end
$scope module ff_1 $end
$var reg 1 4 t $end
$var reg 1 5 en $end
$var reg 1 6 rst $end
$var reg 1 7 clk $end
$var reg 1 8 q $end
$var reg 1 9 q_pres $end
$var reg 1 : q_next $end
$upscope $end
$scope module ff_2 $end
$var reg 1 ; t $end
$var reg 1 < en $end
$var reg 1 = rst $end
$var reg 1 > clk $end
$var reg 1 ? q $end
$var reg 1 @ q_pres $end
$var reg 1 A q_next $end
$upscope $end
$scope module ff_3 $end
$var reg 1 B t $end
$var reg 1 C en $end
$var reg 1 D rst $end
$var reg 1 E clk $end
$var reg 1 F q $end
$var reg 1 G q_pres $end
$var reg 1 H q_next $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
1#
b000 $
0%
0&
1'
b000 (
0)
0*
0+
0,
1-
0.
0/
00
b00000000000000000000 1
b00000000000000000001 2
03
14
15
16
07
08
09
1:
0;
1<
1=
0>
0?
0@
0A
0B
1C
1D
0E
0F
0G
0H
#5000000
1!
0#
1%
0'
0-
1.
06
0=
0D
#10000000
0!
1"
0%
1&
0.
1/
#15000000
1!
1%
1.
b00000000000000000001 1
b00000000000000000010 2
#20000000
0!
0"
0%
0&
0.
0/
#25000000
1!
1%
1.
b00000000000000000010 1
b00000000000000000011 2
#30000000
0!
1"
0%
1&
0.
1/
#35000000
1!
1%
1.
b00000000000000000011 1
b00000000000000000100 2
#40000000
0!
0"
0%
0&
0.
0/
#45000000
1!
1%
1.
b00000000000000000100 1
b00000000000000000101 2
#50000000
0!
1"
0%
1&
0.
1/
#55000000
1!
1%
1.
b00000000000000000101 1
b00000000000000000110 2
#60000000
0!
0"
0%
0&
0.
0/
#65000000
1!
1%
1.
b00000000000000000110 1
b00000000000000000111 2
#70000000
0!
1"
0%
1&
0.
1/
#75000000
1!
1%
1.
b00000000000000000111 1
b00000000000000001000 2
#80000000
0!
0"
0%
0&
0.
0/
#85000000
1!
1%
1.
b00000000000000001000 1
b00000000000000001001 2
#90000000
0!
1"
0%
1&
0.
1/
#95000000
1!
1%
1.
b00000000000000001001 1
b00000000000000001010 2
#100000000
0!
0"
0%
0&
0.
0/
#105000000
1!
1%
1.
b00000000000000001010 1
b00000000000000001011 2
#110000000
0!
1"
0%
1&
0.
1/
#115000000
1!
1%
1.
b00000000000000001011 1
b00000000000000001100 2
#120000000
0!
0"
0%
0&
0.
0/
#125000000
1!
1%
1.
b00000000000000001100 1
b00000000000000001101 2
#130000000
0!
1"
0%
1&
0.
1/
#135000000
1!
1%
1.
b00000000000000001101 1
b00000000000000001110 2
#140000000
0!
0"
0%
0&
0.
0/
#145000000
1!
1%
1.
b00000000000000001110 1
b00000000000000001111 2
#150000000
0!
1"
0%
1&
0.
1/
#155000000
1!
1%
1.
b00000000000000001111 1
b00000000000000010000 2
#160000000
0!
0"
0%
0&
0.
0/
#165000000
1!
1%
1.
b00000000000000010000 1
b00000000000000010001 2
#170000000
0!
1"
0%
1&
0.
1/
#175000000
1!
1%
1.
b00000000000000010001 1
b00000000000000010010 2
#180000000
0!
0"
0%
0&
0.
0/
#185000000
1!
1%
1.
b00000000000000010010 1
b00000000000000010011 2
#190000000
0!
1"
0%
1&
0.
1/
#195000000
1!
1%
1.
b00000000000000010011 1
b00000000000000010100 2
#200000000
0!
0"
0%
0&
0.
0/
#205000000
1!
1%
1.
b00000000000000010100 1
b00000000000000010101 2
#210000000
0!
1"
0%
1&
0.
1/
#215000000
1!
1%
1.
b00000000000000010101 1
b00000000000000010110 2
#220000000
0!
0"
0%
0&
0.
0/
#225000000
1!
1%
1.
b00000000000000010110 1
b00000000000000010111 2
#230000000
0!
1"
0%
1&
0.
1/
#235000000
1!
1%
1.
b00000000000000010111 1
b00000000000000011000 2
#240000000
0!
0"
0%
0&
0.
0/
#245000000
1!
1%
1.
b00000000000000011000 1
b00000000000000011001 2
#250000000
0!
1"
0%
1&
0.
1/
#255000000
1!
1%
1.
b00000000000000011001 1
b00000000000000011010 2
#260000000
0!
0"
0%
0&
0.
0/
#265000000
1!
1%
1.
b00000000000000011010 1
b00000000000000011011 2
#270000000
0!
1"
0%
1&
0.
1/
#275000000
1!
1%
1.
b00000000000000011011 1
b00000000000000011100 2
#280000000
0!
0"
0%
0&
0.
0/
#285000000
1!
1%
1.
b00000000000000011100 1
b00000000000000011101 2
#290000000
0!
1"
0%
1&
0.
1/
#295000000
1!
1%
1.
b00000000000000011101 1
b00000000000000011110 2
