-- VHDL 8 bit processor Project
-- Full Adder (decomposed)
-- James Hicks Sept 21 2023

